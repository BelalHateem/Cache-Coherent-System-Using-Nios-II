-- top.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity top is
	port (
		clk_clk                             : in    std_logic                     := '0';             --                          clk.clk
		reset_reset                         : in    std_logic                     := '0';             --                        reset.reset
		sdram_clk_clk                       : out   std_logic;                                        --                    sdram_clk.clk
		sdram_wire_addr                     : out   std_logic_vector(12 downto 0);                    --                   sdram_wire.addr
		sdram_wire_ba                       : out   std_logic_vector(1 downto 0);                     --                             .ba
		sdram_wire_cas_n                    : out   std_logic;                                        --                             .cas_n
		sdram_wire_cke                      : out   std_logic;                                        --                             .cke
		sdram_wire_cs_n                     : out   std_logic;                                        --                             .cs_n
		sdram_wire_dq                       : inout std_logic_vector(31 downto 0) := (others => '0'); --                             .dq
		sdram_wire_dqm                      : out   std_logic_vector(3 downto 0);                     --                             .dqm
		sdram_wire_ras_n                    : out   std_logic;                                        --                             .ras_n
		sdram_wire_we_n                     : out   std_logic;                                        --                             .we_n
		switches_external_connection_export : in    std_logic_vector(7 downto 0)  := (others => '0')  -- switches_external_connection.export
	);
end entity top;

architecture rtl of top is
	component top_cpu_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component top_cpu_0;

	component top_cpu_1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component top_cpu_1;

	component top_jtag_uart0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component top_jtag_uart0;

	component top_mutex is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component top_mutex;

	component top_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component top_sdram;

	component top_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component top_switches;

	component top_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component top_sys_sdram_pll_0;

	component top_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component top_sysid_qsys;

	component top_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component top_timer_0;

	component top_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                  : in  std_logic                     := 'X';             -- clk
			cpu_0_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			jtag_uart0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart1_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_0_data_master_address                    : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_0_data_master_waitrequest                : out std_logic;                                        -- waitrequest
			cpu_0_data_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_0_data_master_read                       : in  std_logic                     := 'X';             -- read
			cpu_0_data_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_data_master_readdatavalid              : out std_logic;                                        -- readdatavalid
			cpu_0_data_master_write                      : in  std_logic                     := 'X';             -- write
			cpu_0_data_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_0_data_master_debugaccess                : in  std_logic                     := 'X';             -- debugaccess
			cpu_0_instruction_master_address             : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_0_instruction_master_waitrequest         : out std_logic;                                        -- waitrequest
			cpu_0_instruction_master_read                : in  std_logic                     := 'X';             -- read
			cpu_0_instruction_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_instruction_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_address                    : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_1_data_master_waitrequest                : out std_logic;                                        -- waitrequest
			cpu_1_data_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_1_data_master_read                       : in  std_logic                     := 'X';             -- read
			cpu_1_data_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_data_master_readdatavalid              : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_write                      : in  std_logic                     := 'X';             -- write
			cpu_1_data_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_1_data_master_debugaccess                : in  std_logic                     := 'X';             -- debugaccess
			cpu_1_instruction_master_address             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_1_instruction_master_waitrequest         : out std_logic;                                        -- waitrequest
			cpu_1_instruction_master_read                : in  std_logic                     := 'X';             -- read
			cpu_1_instruction_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_instruction_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			cpu_0_debug_mem_slave_address                : out std_logic_vector(8 downto 0);                     -- address
			cpu_0_debug_mem_slave_write                  : out std_logic;                                        -- write
			cpu_0_debug_mem_slave_read                   : out std_logic;                                        -- read
			cpu_0_debug_mem_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_0_debug_mem_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_0_debug_mem_slave_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_0_debug_mem_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			cpu_0_debug_mem_slave_debugaccess            : out std_logic;                                        -- debugaccess
			cpu_1_debug_mem_slave_address                : out std_logic_vector(8 downto 0);                     -- address
			cpu_1_debug_mem_slave_write                  : out std_logic;                                        -- write
			cpu_1_debug_mem_slave_read                   : out std_logic;                                        -- read
			cpu_1_debug_mem_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_1_debug_mem_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_1_debug_mem_slave_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_1_debug_mem_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			cpu_1_debug_mem_slave_debugaccess            : out std_logic;                                        -- debugaccess
			jtag_uart0_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart0_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart0_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart0_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart0_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart0_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart0_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			jtag_uart1_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart1_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart1_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart1_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart1_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart1_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart1_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			mutex_s1_address                             : out std_logic_vector(0 downto 0);                     -- address
			mutex_s1_write                               : out std_logic;                                        -- write
			mutex_s1_read                                : out std_logic;                                        -- read
			mutex_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mutex_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			mutex_s1_chipselect                          : out std_logic;                                        -- chipselect
			sdram_s1_address                             : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                               : out std_logic;                                        -- write
			sdram_s1_read                                : out std_logic;                                        -- read
			sdram_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                          : out std_logic;                                        -- chipselect
			switches_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                             : out std_logic;                                        -- write
			timer_0_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                        : out std_logic;                                        -- chipselect
			timer_1_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                             : out std_logic;                                        -- write
			timer_1_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                        : out std_logic                                         -- chipselect
		);
	end component top_mm_interconnect_0;

	component top_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component top_irq_mapper;

	component top_irq_mapper_001 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component top_irq_mapper_001;

	component top_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component top_rst_controller;

	component top_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component top_rst_controller_001;

	signal sys_sdram_pll_0_sys_clk_clk                                    : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [cpu_0:clk, cpu_1:clk, irq_mapper:clk, irq_mapper_001:clk, jtag_uart0:clk, jtag_uart1:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, mutex:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk, sdram:clk, switches:clk, sysid_qsys:clock, timer_0:clk, timer_1:clk]
	signal cpu_0_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_debugaccess                                  : std_logic;                     -- cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	signal cpu_0_data_master_address                                      : std_logic_vector(27 downto 0); -- cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	signal cpu_0_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	signal cpu_0_data_master_read                                         : std_logic;                     -- cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	signal cpu_0_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	signal cpu_0_data_master_write                                        : std_logic;                     -- cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	signal cpu_0_data_master_writedata                                    : std_logic_vector(31 downto 0); -- cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	signal cpu_1_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	signal cpu_1_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	signal cpu_1_data_master_debugaccess                                  : std_logic;                     -- cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	signal cpu_1_data_master_address                                      : std_logic_vector(27 downto 0); -- cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	signal cpu_1_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	signal cpu_1_data_master_read                                         : std_logic;                     -- cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	signal cpu_1_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	signal cpu_1_data_master_write                                        : std_logic;                     -- cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	signal cpu_1_data_master_writedata                                    : std_logic_vector(31 downto 0); -- cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	signal cpu_0_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                               : std_logic_vector(27 downto 0); -- cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	signal cpu_0_instruction_master_read                                  : std_logic;                     -- cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	signal cpu_0_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	signal cpu_1_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	signal cpu_1_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	signal cpu_1_instruction_master_address                               : std_logic_vector(26 downto 0); -- cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	signal cpu_1_instruction_master_read                                  : std_logic;                     -- cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	signal cpu_1_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart0_avalon_jtag_slave_chipselect -> jtag_uart0:av_chipselect
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart0:av_readdata -> mm_interconnect_0:jtag_uart0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart0:av_waitrequest -> mm_interconnect_0:jtag_uart0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart0_avalon_jtag_slave_address -> jtag_uart0:av_address
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart0_avalon_jtag_slave_writedata -> jtag_uart0:av_writedata
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata            : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest            : std_logic;                     -- cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_0_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	signal mm_interconnect_0_cpu_0_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_0_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	signal mm_interconnect_0_cpu_0_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                          : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_mutex_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:mutex_s1_chipselect -> mutex:chipselect
	signal mm_interconnect_0_mutex_s1_readdata                            : std_logic_vector(31 downto 0); -- mutex:data_to_cpu -> mm_interconnect_0:mutex_s1_readdata
	signal mm_interconnect_0_mutex_s1_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mutex_s1_address -> mutex:address
	signal mm_interconnect_0_mutex_s1_read                                : std_logic;                     -- mm_interconnect_0:mutex_s1_read -> mutex:read
	signal mm_interconnect_0_mutex_s1_write                               : std_logic;                     -- mm_interconnect_0:mutex_s1_write -> mutex:write
	signal mm_interconnect_0_mutex_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:mutex_s1_writedata -> mutex:data_from_cpu
	signal mm_interconnect_0_switches_s1_readdata                         : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_sdram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                            : std_logic_vector(31 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                         : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                             : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                       : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                               : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_cpu_1_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest            : std_logic;                     -- cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_1_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	signal mm_interconnect_0_cpu_1_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_1_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	signal mm_interconnect_0_cpu_1_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart1_avalon_jtag_slave_chipselect -> jtag_uart1:av_chipselect
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart1:av_readdata -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart1:av_waitrequest -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart1_avalon_jtag_slave_address -> jtag_uart1:av_address
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart1_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart1_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart1_avalon_jtag_slave_writedata -> jtag_uart1:av_writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                          : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                             : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                       : std_logic;                     -- jtag_uart0:av_irq -> irq_mapper:receiver1_irq
	signal cpu_0_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_0:irq
	signal irq_mapper_001_receiver0_irq                                   : std_logic;                     -- timer_1:irq -> irq_mapper_001:receiver0_irq
	signal irq_mapper_001_receiver1_irq                                   : std_logic;                     -- jtag_uart1:av_irq -> irq_mapper_001:receiver1_irq
	signal cpu_1_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> cpu_1:irq
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                             : std_logic;                     -- rst_controller:reset_req -> [cpu_0:reset_req, cpu_1:reset_req, rst_translator:reset_req_in]
	signal cpu_0_debug_reset_request_reset                                : std_logic;                     -- cpu_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal cpu_1_debug_reset_request_reset                                : std_logic;                     -- cpu_1:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in0]
	signal sys_sdram_pll_0_reset_source_reset                             : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in2, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                             : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:jtag_uart1_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read:inv -> jtag_uart0:av_read_n
	signal mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write:inv -> jtag_uart0:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read:inv -> jtag_uart1:av_read_n
	signal mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write:inv -> jtag_uart1:av_write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu_0:reset_n, cpu_1:reset_n, mutex:reset_n, sdram:reset_n, switches:reset_n, sysid_qsys:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart0:rst_n, timer_0:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [jtag_uart1:rst_n, timer_1:reset_n]

begin

	cpu_0 : component top_cpu_0
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                         --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_0_data_master_read,                              --                          .read
			d_readdata                          => cpu_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_0_data_master_write,                             --                          .write
			d_writedata                         => cpu_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_1 : component top_cpu_1
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                         --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_1_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_1_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_1_data_master_read,                              --                          .read
			d_readdata                          => cpu_1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_1_data_master_write,                             --                          .write
			d_writedata                         => cpu_1_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_1_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_1_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	jtag_uart0 : component top_jtag_uart0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                    --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                        --               irq.irq
		);

	jtag_uart1 : component top_jtag_uart0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                    --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver1_irq                                    --               irq.irq
		);

	mutex : component top_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv, -- reset.reset_n
			clk           => sys_sdram_pll_0_sys_clk_clk,              --   clk.clk
			chipselect    => mm_interconnect_0_mutex_s1_chipselect,    --    s1.chipselect
			data_from_cpu => mm_interconnect_0_mutex_s1_writedata,     --      .writedata
			read          => mm_interconnect_0_mutex_s1_read,          --      .read
			write         => mm_interconnect_0_mutex_s1_write,         --      .write
			data_to_cpu   => mm_interconnect_0_mutex_s1_readdata,      --      .readdata
			address       => mm_interconnect_0_mutex_s1_address(0)     --      .address
		);

	sdram : component top_sdram
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                     --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	switches : component top_switches
		port map (
			clk      => sys_sdram_pll_0_sys_clk_clk,              --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_external_connection_export       -- external_connection.export
		);

	sys_sdram_pll_0 : component top_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => reset_reset,                        --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	sysid_qsys : component top_sysid_qsys
		port map (
			clock    => sys_sdram_pll_0_sys_clk_clk,                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer_0 : component top_timer_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                      --   irq.irq
		);

	timer_1 : component top_timer_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_001_receiver0_irq                  --   irq.irq
		);

	mm_interconnect_0 : component top_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                  => sys_sdram_pll_0_sys_clk_clk,                                --                sys_sdram_pll_0_sys_clk.clk
			cpu_0_reset_reset_bridge_in_reset_reset      => rst_controller_reset_out_reset,                             --      cpu_0_reset_reset_bridge_in_reset.reset
			jtag_uart0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                         -- jtag_uart0_reset_reset_bridge_in_reset.reset
			jtag_uart1_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                         -- jtag_uart1_reset_reset_bridge_in_reset.reset
			cpu_0_data_master_address                    => cpu_0_data_master_address,                                  --                      cpu_0_data_master.address
			cpu_0_data_master_waitrequest                => cpu_0_data_master_waitrequest,                              --                                       .waitrequest
			cpu_0_data_master_byteenable                 => cpu_0_data_master_byteenable,                               --                                       .byteenable
			cpu_0_data_master_read                       => cpu_0_data_master_read,                                     --                                       .read
			cpu_0_data_master_readdata                   => cpu_0_data_master_readdata,                                 --                                       .readdata
			cpu_0_data_master_readdatavalid              => cpu_0_data_master_readdatavalid,                            --                                       .readdatavalid
			cpu_0_data_master_write                      => cpu_0_data_master_write,                                    --                                       .write
			cpu_0_data_master_writedata                  => cpu_0_data_master_writedata,                                --                                       .writedata
			cpu_0_data_master_debugaccess                => cpu_0_data_master_debugaccess,                              --                                       .debugaccess
			cpu_0_instruction_master_address             => cpu_0_instruction_master_address,                           --               cpu_0_instruction_master.address
			cpu_0_instruction_master_waitrequest         => cpu_0_instruction_master_waitrequest,                       --                                       .waitrequest
			cpu_0_instruction_master_read                => cpu_0_instruction_master_read,                              --                                       .read
			cpu_0_instruction_master_readdata            => cpu_0_instruction_master_readdata,                          --                                       .readdata
			cpu_0_instruction_master_readdatavalid       => cpu_0_instruction_master_readdatavalid,                     --                                       .readdatavalid
			cpu_1_data_master_address                    => cpu_1_data_master_address,                                  --                      cpu_1_data_master.address
			cpu_1_data_master_waitrequest                => cpu_1_data_master_waitrequest,                              --                                       .waitrequest
			cpu_1_data_master_byteenable                 => cpu_1_data_master_byteenable,                               --                                       .byteenable
			cpu_1_data_master_read                       => cpu_1_data_master_read,                                     --                                       .read
			cpu_1_data_master_readdata                   => cpu_1_data_master_readdata,                                 --                                       .readdata
			cpu_1_data_master_readdatavalid              => cpu_1_data_master_readdatavalid,                            --                                       .readdatavalid
			cpu_1_data_master_write                      => cpu_1_data_master_write,                                    --                                       .write
			cpu_1_data_master_writedata                  => cpu_1_data_master_writedata,                                --                                       .writedata
			cpu_1_data_master_debugaccess                => cpu_1_data_master_debugaccess,                              --                                       .debugaccess
			cpu_1_instruction_master_address             => cpu_1_instruction_master_address,                           --               cpu_1_instruction_master.address
			cpu_1_instruction_master_waitrequest         => cpu_1_instruction_master_waitrequest,                       --                                       .waitrequest
			cpu_1_instruction_master_read                => cpu_1_instruction_master_read,                              --                                       .read
			cpu_1_instruction_master_readdata            => cpu_1_instruction_master_readdata,                          --                                       .readdata
			cpu_1_instruction_master_readdatavalid       => cpu_1_instruction_master_readdatavalid,                     --                                       .readdatavalid
			cpu_0_debug_mem_slave_address                => mm_interconnect_0_cpu_0_debug_mem_slave_address,            --                  cpu_0_debug_mem_slave.address
			cpu_0_debug_mem_slave_write                  => mm_interconnect_0_cpu_0_debug_mem_slave_write,              --                                       .write
			cpu_0_debug_mem_slave_read                   => mm_interconnect_0_cpu_0_debug_mem_slave_read,               --                                       .read
			cpu_0_debug_mem_slave_readdata               => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,           --                                       .readdata
			cpu_0_debug_mem_slave_writedata              => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,          --                                       .writedata
			cpu_0_debug_mem_slave_byteenable             => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,         --                                       .byteenable
			cpu_0_debug_mem_slave_waitrequest            => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest,        --                                       .waitrequest
			cpu_0_debug_mem_slave_debugaccess            => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess,        --                                       .debugaccess
			cpu_1_debug_mem_slave_address                => mm_interconnect_0_cpu_1_debug_mem_slave_address,            --                  cpu_1_debug_mem_slave.address
			cpu_1_debug_mem_slave_write                  => mm_interconnect_0_cpu_1_debug_mem_slave_write,              --                                       .write
			cpu_1_debug_mem_slave_read                   => mm_interconnect_0_cpu_1_debug_mem_slave_read,               --                                       .read
			cpu_1_debug_mem_slave_readdata               => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,           --                                       .readdata
			cpu_1_debug_mem_slave_writedata              => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,          --                                       .writedata
			cpu_1_debug_mem_slave_byteenable             => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,         --                                       .byteenable
			cpu_1_debug_mem_slave_waitrequest            => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest,        --                                       .waitrequest
			cpu_1_debug_mem_slave_debugaccess            => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess,        --                                       .debugaccess
			jtag_uart0_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address,     --           jtag_uart0_avalon_jtag_slave.address
			jtag_uart0_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write,       --                                       .write
			jtag_uart0_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read,        --                                       .read
			jtag_uart0_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata,    --                                       .readdata
			jtag_uart0_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata,   --                                       .writedata
			jtag_uart0_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest, --                                       .waitrequest
			jtag_uart0_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect,  --                                       .chipselect
			jtag_uart1_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address,     --           jtag_uart1_avalon_jtag_slave.address
			jtag_uart1_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write,       --                                       .write
			jtag_uart1_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read,        --                                       .read
			jtag_uart1_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata,    --                                       .readdata
			jtag_uart1_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata,   --                                       .writedata
			jtag_uart1_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest, --                                       .waitrequest
			jtag_uart1_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect,  --                                       .chipselect
			mutex_s1_address                             => mm_interconnect_0_mutex_s1_address,                         --                               mutex_s1.address
			mutex_s1_write                               => mm_interconnect_0_mutex_s1_write,                           --                                       .write
			mutex_s1_read                                => mm_interconnect_0_mutex_s1_read,                            --                                       .read
			mutex_s1_readdata                            => mm_interconnect_0_mutex_s1_readdata,                        --                                       .readdata
			mutex_s1_writedata                           => mm_interconnect_0_mutex_s1_writedata,                       --                                       .writedata
			mutex_s1_chipselect                          => mm_interconnect_0_mutex_s1_chipselect,                      --                                       .chipselect
			sdram_s1_address                             => mm_interconnect_0_sdram_s1_address,                         --                               sdram_s1.address
			sdram_s1_write                               => mm_interconnect_0_sdram_s1_write,                           --                                       .write
			sdram_s1_read                                => mm_interconnect_0_sdram_s1_read,                            --                                       .read
			sdram_s1_readdata                            => mm_interconnect_0_sdram_s1_readdata,                        --                                       .readdata
			sdram_s1_writedata                           => mm_interconnect_0_sdram_s1_writedata,                       --                                       .writedata
			sdram_s1_byteenable                          => mm_interconnect_0_sdram_s1_byteenable,                      --                                       .byteenable
			sdram_s1_readdatavalid                       => mm_interconnect_0_sdram_s1_readdatavalid,                   --                                       .readdatavalid
			sdram_s1_waitrequest                         => mm_interconnect_0_sdram_s1_waitrequest,                     --                                       .waitrequest
			sdram_s1_chipselect                          => mm_interconnect_0_sdram_s1_chipselect,                      --                                       .chipselect
			switches_s1_address                          => mm_interconnect_0_switches_s1_address,                      --                            switches_s1.address
			switches_s1_readdata                         => mm_interconnect_0_switches_s1_readdata,                     --                                       .readdata
			sysid_qsys_control_slave_address             => mm_interconnect_0_sysid_qsys_control_slave_address,         --               sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata            => mm_interconnect_0_sysid_qsys_control_slave_readdata,        --                                       .readdata
			timer_0_s1_address                           => mm_interconnect_0_timer_0_s1_address,                       --                             timer_0_s1.address
			timer_0_s1_write                             => mm_interconnect_0_timer_0_s1_write,                         --                                       .write
			timer_0_s1_readdata                          => mm_interconnect_0_timer_0_s1_readdata,                      --                                       .readdata
			timer_0_s1_writedata                         => mm_interconnect_0_timer_0_s1_writedata,                     --                                       .writedata
			timer_0_s1_chipselect                        => mm_interconnect_0_timer_0_s1_chipselect,                    --                                       .chipselect
			timer_1_s1_address                           => mm_interconnect_0_timer_1_s1_address,                       --                             timer_1_s1.address
			timer_1_s1_write                             => mm_interconnect_0_timer_1_s1_write,                         --                                       .write
			timer_1_s1_readdata                          => mm_interconnect_0_timer_1_s1_readdata,                      --                                       .readdata
			timer_1_s1_writedata                         => mm_interconnect_0_timer_1_s1_writedata,                     --                                       .writedata
			timer_1_s1_chipselect                        => mm_interconnect_0_timer_1_s1_chipselect                     --                                       .chipselect
		);

	irq_mapper : component top_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_0_irq_irq                   --    sender.irq
		);

	irq_mapper_001 : component top_irq_mapper_001
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,   -- receiver0.irq
			receiver1_irq => irq_mapper_001_receiver1_irq,   -- receiver1.irq
			sender_irq    => cpu_1_irq_irq                   --    sender.irq
		);

	rst_controller : component top_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_0_debug_reset_request_reset,    -- reset_in0.reset
			reset_in1      => cpu_1_debug_reset_request_reset,    -- reset_in1.reset
			reset_in2      => sys_sdram_pll_0_reset_source_reset, -- reset_in2.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component top_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_0_debug_reset_request_reset,    -- reset_in0.reset
			reset_in1      => sys_sdram_pll_0_reset_source_reset, -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component top_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_1_debug_reset_request_reset,    -- reset_in0.reset
			reset_in1      => sys_sdram_pll_0_reset_source_reset, -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of top
